`timescale 1ns / 1ps
module tb();

////////////////////////
// Local declarations //
////////////////////////

    parameter              PERIOD     = 83.3;
    parameter              LENGTH     = 63;             //code lenght for checks   
    parameter              POLY_LEN   = $clog2(LENGTH); //polynom lenght 
    parameter              HOLD_PARAM = 3;

    logic                  clkin;                       //clocking
    logic                  rstn;                        //reset
   
    logic [POLY_LEN-1:0]   code1;                //phase signals

    logic [LENGTH-1:0]     final_gold_code;             //the register that serves to check the final Gold code       

    logic                  code_gold;                   //1 bit of Gold code
    logic [LENGTH-1:0]     ref_code;                    //Reference code for comparison

    integer                shift_state;
    integer                shift;
    integer                hold;
    
    logic [LENGTH-1:0] table_gold[0:LENGTH];            //Table of values 
    axistream_if        axis(clkin);       

/////////////////
// Connections //
/////////////////

    Gold_gen gold_gen(
        .clkin(clkin),
        .rstn(rstn), 
        .code_gold(code_gold),
        .strobe_sig_o(),
        .s_axis(axis)
    );

////////////////
// Test bench //
///////////////

//clk simulation
    initial forever begin
          #(PERIOD/2) clkin = 1'b1;
          #(PERIOD/2) clkin = 1'b0;
    end

//Results saving block and start values
    initial begin
    shift_state <= 0;
        rstn <= 0;
        hold <= HOLD_PARAM - 1;
        axis.tvalid <= 1;
        #100;
        rstn <= 1;
        #10
        code1 <= 6'b000000;
        axis.tdata <= 6'b000000;
    
    table_gold = '{63'b000000110011000000001101010101110101000000101010011101101000001, 63'b111111100100000110010000110101001001100101111001001101001010111, 63'b000001001010001010101011110100110000101111011111101100001111010, 63'b111100010110010011011101110111000010111010010010101110000100001, 
    63'b000110101110100000110001110000100110010000001000101010010010110, 63'b110011011111000111101001111111101111000100111100100010111111001, 63'b011000111100001001011001100001111101101101010100110011100100110, 63'b001111111010010100111001011101011000111110000100010001010011001, 63'b100001110110101111111000100100010010011000100101010100111100111, 
    63'b111101101111011001111011010110000111010101100111011111100011010, 63'b000101011100110101111100110010101101001111100011001001011100000, 63'b110100111011101101110011111011111001111011101011100100100010101, 63'b010111110101011101101101101001010000010011111010111111011111110, 63'b010001101000111101010001001100000011000011011000001000100101001, 
    63'b011101010011111100101000000110100101100010011101100111010000111, 63'b000100100101111111011010010011101000100000010110111000111011011, 63'b110111001001111000111110111001110010100100000000000111101100011, 63'b010000010001110111110111101101000110101100101101111001000010010, 63'b011110100001101001100101000100101110111101110110000100011110001, 
    63'b000011000001010101000000010111111110011111000001111110100110111, 63'b111000000000101100001010110001011111011010101110001011010111011, 63'b001110000011011110011111111100011101010001110001100000110100010, 63'b100010000100111010110101100110011001000111001110110111110010001, 63'b111010001011110011100001010010010001101010110000011001111110110, 
    63'b001010010101100001001000111010000000110001001101000101100111000, 63'b101010101001000100011011101010100010000110110111111101010100101, 63'b101011010000001110111101001011100111101001000010001100110011110, 63'b101000100010011011110000001001101100110110101001101111111101000, 63'b101111000110110001101010001101111010001001111110101001100000100, 
    63'b100000001111100101011110000101010111110111010000100101011011100, 63'b111110011101001100110110010100001100001010001100111100101101100, 63'b000010111000011111100110110110111011110000110100001111000001100, 63'b111011110010111001000111110011010100000101000101101000011001101, 63'b001001100111110100000101111000001011101110100110100110101001110, 
    63'b101101001101101110000001101110110100111001100000111011001001001, 63'b100100011001011010001001000011001010010111101100000000001000110, 63'b110110110000110010011000011000110111001011110101110110001011000, 63'b010011100011100010111010101111001101110011000110011010001100100, 63'b011001000101000011111111000000111000000010100001000010000011101, 
    63'b001100001000000001110100011111010011100001101111110010011101111, 63'b100110010010000101100010100000000100100111110010010010100001011, 63'b110010100110001101001111011110101010101011001001010011011000010, 63'b011011001110011100010100100011110110110010111111010000101010000, 63'b001000011110111110100011011001001110000001010011010111001110101, 
    63'b101110111111111011001100101100111111100110001011011000000111111, 63'b100011111101110000010011000111011100101000111011000110010101010, 63'b111001111001100110101100010000011010110101011011111010110000000, 63'b001101110001001011010010111110010110001110011010000011111010100, 63'b100101100000010000101111100010001111111000011001110001101111101, 
    63'b110101000010100111010101011010111100010100011110010101000101110, 63'b010100000111001000100000101011011011001100010001011100010001000, 63'b010110001100010111001011001000010101111100001111001110111000101, 63'b010010011010101000011100001110001000011100110011101011101011111, 63'b011010110111010110110010000010110011011101001010100001001101011, 
    63'b001011101100101011101110011011000101011110111000110100000000011, 63'b101001011011010001010110101000101001011001011100011110011010011, 63'b101100110100100100100111001111110001010110010101001010101110010, 63'b100111101011001111000100000001000001001000000111100011000110000, 63'b110001010100011000000010011100100001110100100010110000010110100, 
    63'b011100101010110110001110100111100000001101101000010110110111100, 63'b000111010111101010010111010001100011111111111101011011110101101, 63'b110000101101010010100100111101100100011011010111000001110001111, 63'b011111011000100011000011100101101011010010000011110101111001010, 63'b000000110011000000001101010101110101000000101010011101101000001};
         
        forever begin
                @(posedge clkin);
                while (!axis.tready) begin
                   @(posedge clkin);
                end
                
                shift = shift_state;
                ref_code = table_gold[shift];
                
                repeat ((LENGTH+2) * HOLD_PARAM) begin         
                    if(hold != 0) begin
                        hold <= hold - 1;
                    end else begin 
                        final_gold_code <= {final_gold_code[LENGTH-2:0], code_gold};
                        hold <= HOLD_PARAM - 1;                  
                    end
                    @(posedge clkin);
                end
                    
                if(final_gold_code == ref_code) begin
                    $display("Shift %0d is correct!", shift);
                end else begin
                    $display("Shift %0d is incorrect!", shift);
                end  
            end
        end

//code2 initial change block
        initial begin
            forever begin 
            
              while (!axis.tready) begin
                    @(posedge clkin);
              end
              
              repeat ((LENGTH-2) * HOLD_PARAM) @(posedge clkin);
              
              shift_state = $urandom_range(0,LENGTH);
              axis.tdata = shift_state;
              
            end 
        end

endmodule
